// uINST_LIST

parameter iBUSA_H = 33,
parameter iBUSA_L = 28,
parameter iBUSB_H = 27,
parameter iBUSB_L = 22,
parameter iBUSC_H = 21,
parameter iBUSC_L = 16,
parameter iALUC_H = 15,
parameter iALUC_L = 12,
parameter iSH_H   = 11,
parameter iSH_L   = 10,
parameter iKMX    = 9,
parameter iT_H    = 8,
parameter iT_L    = 2,
parameter iM_H    = 1,
parameter iM_L    = 0,
//                      AAAAAA_BBBBBB_CCCCCC_ALUC_SH_K_TTTTTTT_MM
// X0000                AAAAAA_BBBBBB_CCCCCC_ALUC_SH_K_TTTTTTT_MM
parameter BSR_u   = 34'b111111_111111_111111_0000_00_0_1000000_00,
parameter MOVMw_u = 34'b111111_111111_111111_0000_00_0_0000001_10,
parameter MOVwM_u = 34'b111111_111111_111110_0000_00_0_0000010_01,

parameter MOVwK_u = 34'b111111_111111_111101_0000_00_1_0000010_00,
parameter ANDwK_u = 34'b111111_111101_111101_0111_00_1_0000011_00,
parameter ORwK_u  = 34'b111111_111101_111101_0110_00_1_0000011_00,
parameter ADDwK_u = 34'b111111_111101_111101_0101_00_1_0110011_00,

parameter RET_u   = 34'b111111_111111_111111_0000_00_0_1000000_00,

parameter JMP_u   = 34'b111111_111111_111111_0000_00_0_1000000_00,
parameter JZE_u   = 34'b111111_111111_111111_0000_00_0_1000001_00,
parameter JNE_u   = 34'b111111_111111_111111_0000_00_0_1000001_00,
parameter JCY_u   = 34'b111111_111111_111111_0000_00_0_1010000_00,

// 0X000                AAAAAA_BBBBBB_CCCCCC_ALUC_SH_K_TTTTTTT_MM
parameter MOVij_u = 34'b111111_111111_111111_0000_00_0_0001100_00,
parameter ADDij_u = 34'b111111_111101_111111_0101_00_0_0111101_00,

// 00X00                AAAAAA_BBBBBB_CCCCCC_ALUC_SH_K_TTTTTTT_MM
parameter MOViw_u = 34'b111111_111101_111111_0001_00_0_0001001_00,

parameter MOVwj_u = 34'b111111_111111_111101_0000_00_0_0000110_00,
parameter ANDwj_u = 34'b111111_111101_111101_0111_00_0_0000111_00,
parameter ORwj_u  = 34'b111111_111101_111101_0110_00_0_0000111_00,
parameter ADDwj_u = 34'b111111_111101_111101_0101_00_0_0110111_00,

parameter CPLi_u  = 34'b111111_111111_111111_0010_00_0_0001100_00,
parameter SHLi_u  = 34'b111111_111111_111111_0000_01_0_0001100_00,
parameter SHRi_u  = 34'b111111_111111_111111_0000_10_0_0001100_00,
parameter ASRi_u  = 34'b111111_111111_111111_0000_11_0_0001100_00,

parameter INCi_u  = 34'b111111_111111_111111_1101_00_0_0101100_00,
parameter DECi_u  = 34'b111111_111111_111111_1110_00_0_0101100_00,

// 000X0                AAAAAA_BBBBBB_CCCCCC_ALUC_SH_K_TTTTTTT_MM
parameter CLC_u   = 34'b111111_111111_111111_1011_00_0_0100000_00,
parameter SEC_u   = 34'b111111_111111_111111_1100_00_0_0100000_00,

parameter CPLw_u  = 34'b111111_111101_111101_0011_00_0_0000011_00,
parameter SHLw_u  = 34'b111111_111101_111101_0001_01_0_0000011_00,
parameter SHRw_u  = 34'b111111_111101_111101_0001_10_0_0000011_00,
parameter ASRw_u  = 34'b111111_111101_111101_0001_11_0_0000011_00,

parameter INCw_u  = 34'b111101_111111_111101_1101_00_0_0100011_00,
parameter DECw_u  = 34'b111101_111111_111101_1110_00_0_0100011_00,

parameter NOP_u   = 34'b111111_111111_111111_0000_00_0_0000000_00
